module main

import lib.lex
import log

fn main() {
	lex.add(1, 1)
}

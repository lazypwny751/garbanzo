module lex

pub fn add(a int, b int) {
	println(a + b)
}
